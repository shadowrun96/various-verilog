module hello(A,B);

	input A;
	output B;

	assign B = A;

endmodule
